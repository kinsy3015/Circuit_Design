module m_can_tb();
endmodule