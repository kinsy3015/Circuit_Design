module behavior_tb2();
endmodule